entity minha_entidade is 
    port(signal-nomes: mode signal type;//"signal-name" nome da porta
    signal-names: mode signal type;//"mode" in,out,inout
    signal-names: mode signal type);
end minha_entidade;
          
